*LM111
*Sngl Differential Comp pkg:DIP8 2,3,8,4,7,1
*
* Connections:
*             Non-Inverting Input
*             |   Inverting Input
*             |   |   Positive Power Supply
*             |   |   |   Negative power Supply
*             |   |   |   |   Out+
*             |   |   |   |   |   Out-
*             |   |   |   |   |   |
.SUBCKT LM111 1   2   3   4   5   6
F1  9  3 V1 1
IEE 3  7 DC 100E-6
VI1 21  1 DC .45
VI2 22  2 DC .45
Q1  9 21  7 QIN
Q2  8 22  7 QIN
Q3  9  8  4 QMO
Q4  8  8  4 QMI
.MODEL QIN PNP(IS=800E-18 BF=833.3)
.MODEL QMI NPN(IS=800E-18 BF=1002)
.MODEL QMO NPN(IS=800E-18 BF=1000 CJC=1E-15 TR=118.8E-9)
E1 10  6  9  4  1
V1 10 11 DC 0
Q5  5 11  6 QOC
.MODEL QOC NPN(IS=800E-18 BF=34.49E3 CJC=1E-15 TF=364.6E-12 TR=79.34E-9)
DP  4  3 DX
RP  3  4 6.122E3
.MODEL DX D(IS=800E-18 RS=1)
.ENDS LM111