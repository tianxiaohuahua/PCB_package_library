* TLC3702 VOLTAGE COMPARATOR "MACROMODEL" SUBCIRCUIT
* CREATED USING PARTS VERSION 4.03 ON 03/14/90 AT 10:09
* REV (N/A)
* NOTE: COMPONENTS ADDED TO SIMULATE ACTIVE PULL-UP
* CONNECTIONS:   NON-INVERTING INPUT
*                | INVERTING INPUT
*                | | POSITIVE POWER SUPPLY
*                | | | NEGATIVE POWER SUPPLY
*                | | | | OUTPUT
*                | | | | |
.SUBCKT TLC3702  1 2 3 4 5
  F1    9  3 V1 1

  *THESE COMPONENTS ADDED TO SIMULATE ACTIVE PULL-UP
  *FOUT 30 5 POLY(1) (V1) 4E-3 -40
    BFOUT 30 5 I=4E-3-40*I(V1)
  *EO1 30 0 POLY(1) (3,0) -.75 1
    BEO1 30 0 V=-0.75+1*v(3,0)
    DO1 5  30  DX

  IEE   3  7 DC 100.0E-6
  VI1  21  1 DC .75
  VI2  22  2 DC .75
  Q1    9 21  7 QIN
  Q2    8 22  7 QIN
  Q3    9  8  4 QMO
  Q4    8  8  4 QMI
.MODEL QIN PNP(IS=800.0E-18 BF=10.00E6)
.MODEL QMI NPN(IS=800.0E-18 BF=1002)
.MODEL QMO NPN(IS=800.0E-18 BF=1000 CJC=1E-15 TR=807.4E-9)
  E1   10  4  9  4  1
  V1   10 11 DC 0
  Q5    5 11  4 QOC
.MODEL QOC NPN(IS=800.0E-18 BF=1.810E3 CJC=1E-15 TF=1.357E-9 TR=1.129E-6)
  DP    4  3 DX
  RP 3  4 -70E3
.MODEL DX  D(IS=800.0E-18)
.ENDS TLC3702